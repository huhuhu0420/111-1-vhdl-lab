library ieee;
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.lab8_package.all;

entity lab8 is
	generic (N: integer:=8);
    port (
		clk: in std_logic;
		data: in std_logic_vector(7 downto 0);
		opcode: in std_logic_vector(3 downto 0);
		rs, rt: in std_logic_vector(1 downto 0);
		hex0: out std_logic_vector(6 downto 0);
		hex1: out std_logic_vector(6 downto 0);
		hex2: out std_logic_vector(6 downto 0);
		hex3: out std_logic_vector(6 downto 0);
		hex4: out std_logic_vector(6 downto 0);
		hex5: out std_logic_vector(6 downto 0)
    );
end lab8;

architecture dosth of lab8 is
	TYPE state_type is (load, move, add, andand, sub1, sub2, slt, done);
	TYPE r_type is array (3 downto 0) of std_logic_vector(7 downto 0);
	signal state : state_type := done;
	signal counter : std_logic :='0';
	signal loadCounter: integer := 0;
	signal rsIndex: integer := 0;
	signal rtIndex: integer := 0;
	signal rsOut: std_logic_vector(7 downto 0) := "00000000";
	signal rtOut: std_logic_vector(7 downto 0) := "00000000";
	signal busOut: std_logic_vector(7 downto 0) := "00000000";

begin
	
	process(counter, clk)
	variable r: r_type := (others => (others => '0'));
	begin
		rsIndex <= to_integer(unsigned(rs));
		rtIndex <= to_integer(unsigned(rt));
		busOut <= data;

		if (rising_edge(clk)) then
			if(counter = '1') then
				counter <= '0';
			else 
				counter <= '1';
			end if;
		end if;

		if (rising_edge(counter)) then 
			if state = done then
				case(opcode) is
					when "0000" => state <= load;
					when "0001" => state <= move;
					when "0010" => state <= add;
					when "0011" => state <= andand;
					when "0101" => state <= sub1;
					when "1001" => state <= sub2;
					when "0100" => state <= slt;
					when others => state <= done;
				end case;
			end if;

			case(state) is
				when load =>
					r(rsIndex) := data;
					state <= done;


				when move =>
					r(rsIndex) := r(rtIndex);
					state <= done;

				when add =>
					r(rsIndex) := r(rsIndex) + r(rtIndex);
					state <= done;

				when andand =>
					r(rsIndex) := r(rsIndex) and r(rtIndex);
					state <= done;

				when sub1 =>
					r(rsIndex) := r(rsIndex) - r(rtIndex);
					state <= done;

				when sub2 =>
					r(rsIndex) := r(rtIndex) - r(rsIndex) ;
					state <= done;

				when slt =>
					if r(rsIndex) <r(rtIndex) then
						r(rsIndex) := "00000001";
					else 
						r(rsIndex) := "00000000";
					end if ;
					state <= done;

				when done =>

				when others =>

			end case ;

		end if;
	
	rsOut <= r(rsIndex);
	rtOut <= r(rtIndex);
	busOut <= data;
		
	end process;

	hexRs1: hex port map(rsOut(0), rsOut(1), rsOut(2), rsOut(3), hex2(0), hex2(1), hex2(2), hex2(3), hex2(4), hex2(5), hex2(6));
	hexRs2: hex port map(rsOut(4), rsOut(5), rsOut(6), rsOut(7), hex3(0), hex3(1), hex3(2), hex3(3), hex3(4), hex3(5), hex3(6));
	hexRt1: hex port map(rtOut(0), rtOut(1), rtOut(2), rtOut(3), hex4(0), hex4(1), hex4(2), hex4(3), hex4(4), hex4(5), hex4(6));
	hexRt2: hex port map(rtOut(4), rtOut(5), rtOut(6), rtOut(7), hex5(0), hex5(1), hex5(2), hex5(3), hex5(4), hex5(5), hex5(6));
	hexBus1: hex port map(busOut(0), busOut(1), busOut(2), busOut(3), hex0(0), hex0(1), hex0(2), hex0(3), hex0(4), hex0(5), hex0(6));
	hexBus2: hex port map(busOut(4), busOut(5), busOut(6), busOut(7), hex1(0), hex1(1), hex1(2), hex1(3), hex1(4), hex1(5), hex1(6));

end dosth;